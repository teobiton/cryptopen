`define SPARTAN7