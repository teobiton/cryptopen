`define GENESYSII
// include KINTEX7 specific code (relevant for KC705, GENESYSII,...)
`define KINTEX7